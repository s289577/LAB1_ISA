library verilog;
use verilog.vl_types.all;
entity tb_riscv32i is
end tb_riscv32i;
